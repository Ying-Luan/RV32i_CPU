`timescale 1ns / 1ps

module uart(  // TODO

       );

endmodule
