`timescale 1ns / 1ps

module csr (
           input wire clk,
           input wire rst_n
       );

endmodule
