`timescale 1ns / 1ps

module CSR (
           input wire clk,
           input wire rst_n
       );

endmodule
